library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity po_machine is
    port (
        
    );
end entity po_machine;
